<svg width="50" height="50" viewBox="0 0 100 100" xmlns="http://www.w3.org/2000/svg">
  <title>PortalProje Logo</title>
  <!-- Big navy circle -->
  <circle cx="50" cy="50" r="50" fill="#0a1633" />
  <!-- White "PP" text in center -->
  <text
    x="50%"
    y="55%"
    font-size="40"
    font-weight="bold"
    text-anchor="middle"
    fill="#fff"
    font-family="Arial, sans-serif"
  >
    PP
  </text>
</svg>
